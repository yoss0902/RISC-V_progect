module rnd_rrbn_arb();
